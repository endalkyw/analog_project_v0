.SUBCKT nmos_cm_0 d0 d1 s

* Net:s ----------------


R1 s s:19 2.772
R2 s s:18 0.756
R3 s s:13 1.092
R4 s s:4 3.724
R5 s:4 s:0 32.424
R6 s:4 s:1 3.724
R7 s:4 s:2 0.644
R8 s:2 s:27 2.772
R9 s:2 MN0@2:s 14
R10 s:2 s:26 0.756
R11 s:2 MN0@2:s 14
R12 s:2 s:3 4.368
R13 s:2 MN0@2:s 14
R14 s:3 s:35 2.772
R15 s:3 MN1@2:s 14
R16 s:3 s:34 0.756
R17 s:3 MN1@2:s 14
R18 s:3 s:14 1.092
R19 s:3 MN1@2:s 14
R20 s:34 s:11 1.372
R21 s:34 MN1@2:s 14
R22 s:35 s:36 3.528
R23 s:35 MN1@2:s 14
R24 s:36 s:37 3.528
R25 s:36 MN1@2:s 14
R26 s:37 s:38 3.528
R27 s:37 MN1@2:s 14
R28 s:38 s:39 3.528
R29 s:38 MN1@2:s 14
R30 s:39 s:40 3.528
R31 s:39 MN1@2:s 14
R32 s:40 s:41 3.528
R33 s:40 MN1@2:s 14
R34 s:41 s:12 1.092
R35 s:41 MN1@2:s 14
R36 s:26 s:9 1.372
R37 s:26 MN0@2:s 14
R38 s:27 s:28 3.528
R39 s:27 MN0@2:s 14
R40 s:28 s:29 3.528
R41 s:28 MN0@2:s 14
R42 s:29 s:30 3.528
R43 s:29 MN0@2:s 14
R44 s:30 s:31 3.528
R45 s:30 MN0@2:s 14
R46 s:31 s:32 3.528
R47 s:31 MN0@2:s 14
R48 s:32 s:33 3.528
R49 s:32 MN0@2:s 14
R50 s:33 s:10 1.092
R51 s:33 MN0@2:s 14
R52 s:1 s:19 2.772
R53 s:1 MN0:s 14
R54 s:1 s:18 0.756
R55 s:1 MN0:s 14
R56 s:1 s:13 1.092
R57 s:1 MN0:s 14
R58 s:18 s:7 1.372
R59 s:18 MN0:s 14
R60 s:19 s:20 3.528
R61 s:19 MN0:s 14
R62 s:20 s:21 3.528
R63 s:20 MN0:s 14
R64 s:21 s:22 3.528
R65 s:21 MN0:s 14
R66 s:22 s:23 3.528
R67 s:22 MN0:s 14
R68 s:23 s:24 3.528
R69 s:23 MN0:s 14
R70 s:24 s:25 3.528
R71 s:24 MN0:s 14
R72 s:25 s:8 1.092
R73 s:25 MN0:s 14
R74 s:0 s:15 1.176
R75 s:0 MN0:b 14
R76 s:0 s:16 1.12
R77 s:0 MN0:b 14
R78 s:0 s:17 2.408
R79 s:0 MN0:b 14
R80 s:17 s:6 1.187
R81 s:17 MN0:b 14
R82 s:16 s:5 1.187
R83 s:16 MN0:b 14
R84 MN0:b MN0@2:b 0.01
R85 MN0@2:b MN1:b 0.01
R86 MN1:b MN1@2:b 0.01
R87 MN0@2:s MN1:s 0.01
C1 s:4 0 2.4318000000000003e-13
C2 s:4 0 2.793e-14
C3 s:4 0 4.83e-15
C4 s:2 0 2.0790000000000002e-14
C5 s:2 0 5.67e-15
C6 s:2 0 3.2760000000000004e-14
C7 s:3 0 2.0790000000000002e-14
C8 s:3 0 5.67e-15
C9 s:3 0 8.190000000000001e-15
C10 s:34 0 1.0290000000000001e-14
C11 s:35 0 2.6460000000000002e-14
C12 s:36 0 2.6460000000000002e-14
C13 s:37 0 2.6460000000000002e-14
C14 s:38 0 2.6460000000000002e-14
C15 s:39 0 2.6460000000000002e-14
C16 s:40 0 2.6460000000000002e-14
C17 s:41 0 8.190000000000001e-15
C18 s:26 0 1.0290000000000001e-14
C19 s:27 0 2.6460000000000002e-14
C20 s:28 0 2.6460000000000002e-14
C21 s:29 0 2.6460000000000002e-14
C22 s:30 0 2.6460000000000002e-14
C23 s:31 0 2.6460000000000002e-14
C24 s:32 0 2.6460000000000002e-14
C25 s:33 0 8.190000000000001e-15
C26 s:1 0 2.0790000000000002e-14
C27 s:1 0 5.67e-15
C28 s:1 0 8.190000000000001e-15
C29 s:18 0 1.0290000000000001e-14
C30 s:19 0 2.6460000000000002e-14
C31 s:20 0 2.6460000000000002e-14
C32 s:21 0 2.6460000000000002e-14
C33 s:22 0 2.6460000000000002e-14
C34 s:23 0 2.6460000000000002e-14
C35 s:24 0 2.6460000000000002e-14
C36 s:25 0 8.190000000000001e-15
C37 s:0 0 8.82e-15
C38 s:0 0 8.400000000000001e-15
C39 s:0 0 1.806e-14
C40 s:17 0 8.904000000000007e-15
C41 s:16 0 8.903999999999996e-15


* Net:d0 ----------------


R88 d0 d0:4 0.644
R89 d0 d0:1 0.728
R90 d0:4 d0:5 3.528
R91 d0:4 MN0:d 14
R92 d0:5 d0:6 3.528
R93 d0:5 MN0:d 14
R94 d0:6 d0:7 3.528
R95 d0:6 MN0:d 14
R96 d0:7 d0:8 3.528
R97 d0:7 MN0:d 14
R98 d0:8 d0:9 3.528
R99 d0:8 MN0:d 14
R100 d0:9 d0:10 3.528
R101 d0:9 MN0:d 14
R102 d0:10 d0:11 3.528
R103 d0:10 MN0:d 14
R104 d0:11 d0:0 3.36
R105 d0:11 MN0:d 14
R106 d0:0 d0:2 3.276
R107 d0:0 MN0:g 342
R108 d0:0 MN0@2:g 342
R109 d0:0 MN1:g 342
R110 d0:0 MN1@2:g 342
R111 d0:0 d0:12 0.63
R112 d0:0 MN0:g 342
R113 d0:0 MN0@2:g 342
R114 d0:0 MN1:g 342
R115 d0:0 MN1@2:g 342
R116 d0:12 d0:13 3.528
R117 d0:12 MN0:g 342
R118 d0:12 MN0@2:g 342
R119 d0:12 MN1:g 342
R120 d0:12 MN1@2:g 342
R121 d0:13 d0:3 3.486
R122 d0:13 MN0:g 342
R123 d0:13 MN0@2:g 342
R124 d0:13 MN1:g 342
R125 d0:13 MN1@2:g 342
R126 MN0:d MN0@2:d 0.01
C42 d0:4 0 2.6460000000000002e-14
C43 d0:5 0 2.6460000000000002e-14
C44 d0:6 0 2.6460000000000002e-14
C45 d0:7 0 2.6460000000000002e-14
C46 d0:8 0 2.6460000000000002e-14
C47 d0:9 0 2.6460000000000002e-14
C48 d0:10 0 2.6460000000000002e-14
C49 d0:11 0 2.5200000000000002e-14
C50 d0:0 0 2.457e-14
C51 d0:0 0 4.725e-15
C52 d0:12 0 2.6460000000000002e-14
C53 d0:13 0 2.6145000000000002e-14


* Net:d1 ----------------


R127 d1 d1:5 2.324
R128 d1 d1:1 0.588
R129 d1 d1:3 0.728
R130 d1 d1:4 0.728
R131 d1:4 d1:0 0.728
R132 d1:0 d1:5 2.324
R133 d1:0 d1:1 0.588
R134 d1:0 d1:3 0.728
R135 d1:5 d1:6 3.528
R136 d1:5 MN1:d 14
R137 d1:6 d1:7 3.528
R138 d1:6 MN1:d 14
R139 d1:7 d1:8 3.528
R140 d1:7 MN1:d 14
R141 d1:8 d1:9 3.528
R142 d1:8 MN1:d 14
R143 d1:9 d1:10 3.528
R144 d1:9 MN1:d 14
R145 d1:10 d1:11 3.528
R146 d1:10 MN1:d 14
R147 d1:11 d1:12 3.528
R148 d1:11 MN1:d 14
R149 d1:12 d1:2 1.092
R150 d1:12 MN1:d 14
R151 MN1:d MN1@2:d 0.01
C54 d1:4 0 5.46e-15
C55 d1:0 0 1.743e-14
C56 d1:0 0 4.41e-15
C57 d1:0 0 5.46e-15
C58 d1:5 0 2.6460000000000002e-14
C59 d1:6 0 2.6460000000000002e-14
C60 d1:7 0 2.6460000000000002e-14
C61 d1:8 0 2.6460000000000002e-14
C62 d1:9 0 2.6460000000000002e-14
C63 d1:10 0 2.6460000000000002e-14
C64 d1:11 0 2.6460000000000002e-14
C65 d1:12 0 8.190000000000001e-15


XXMN0 MN0:d MN0:g MN0:s MN0:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=20 nf=1
+ plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=2 par_nf=2 m=1 par=1
+ dtemp=0 l_shape=0 l_shape_s=0 asej=1.188e-14 adej=5.94e-15 psej=2.38e-06
+ pdej=1.08e-06 sca=3.42607 scb=0.000112243 scc=4.33139e-09 lle_sa=3.05e-07
+ lle_sb=7.1e-08 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.695e-06 lle_rxrxb=1.929e-06 lle_rxrxs=1e-06 lle_rxrxn=6.17e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=5.07e-07 lle_ctse=5.07e-07
+ lle_ctnw=2.73e-07 lle_ctsw=2.73e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.252 $Y=0.127
XXMN0@2 MN0@2:d MN0@2:g MN0@2:s MN0@2:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=20
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=2 par_nf=2 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=5.94e-15 adej=5.94e-15 psej=1.08e-06
+ pdej=1.08e-06 sca=3.42607 scb=0.000112243 scc=4.33139e-09 lle_sa=2.27e-07
+ lle_sb=1.49e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.773e-06 lle_rxrxb=1.851e-06 lle_rxrxs=1e-06 lle_rxrxn=2.44079e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=4.29e-07 lle_ctse=4.29e-07
+ lle_ctnw=3.51e-07 lle_ctsw=3.51e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.33 $Y=0.127
XXMN1 MN1:d MN1:g MN1:s MN1:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=20 nf=1
+ plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=2 par_nf=2 m=1 par=1
+ dtemp=0 l_shape=0 l_shape_s=0 asej=5.94e-15 adej=5.94e-15 psej=1.08e-06
+ pdej=1.08e-06 sca=3.42607 scb=0.000112243 scc=4.33139e-09 lle_sa=1.49e-07
+ lle_sb=2.27e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.851e-06 lle_rxrxb=1.773e-06 lle_rxrxs=1e-06 lle_rxrxn=2.44079e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=3.51e-07 lle_ctse=3.51e-07
+ lle_ctnw=4.29e-07 lle_ctsw=4.29e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.408 $Y=0.127
XXMN1@2 MN1@2:d MN1@2:g MN1@2:s MN1@2:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=20
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=2 par_nf=2 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=5.94e-15 adej=1.188e-14
+ psej=1.08e-06 pdej=2.38e-06 sca=3.42607 scb=0.000112243 scc=4.33139e-09
+ lle_sa=7.1e-08 lle_sb=3.05e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06
+ lle_nwn=2e-06 lle_rxrxa=1.929e-06 lle_rxrxb=1.695e-06 lle_rxrxs=1e-06
+ lle_rxrxn=6.17e-07 lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=2.73e-07
+ lle_ctse=2.73e-07 lle_ctnw=5.07e-07 lle_ctsw=5.07e-07 lle_sctne=0 lle_sctnw=0
+ lle_sctse=0 lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.486 $Y=0.127

.ends nmos_cm_0
