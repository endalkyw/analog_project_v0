This is a source file		$must have a title line

.LIB "/project/ssstudents/TAPO_downloads/GF12_V1.0_4.1/12LP/V1.0_4.1/Models/HSPICE/models/12LP_Hspice.lib" TT
.option post = 2
.PARAM wireopt=3 pre_layout_sw=0

.include "../circuits/nmos_cm/nmos_cm_4.sp"
.param vd0_val = 0.8
.param vd1_val = 0.8

xcm d0 d1 0 nmos_cm_4
Vd0 d0 0 DC vd0_val
Vd1 d10 0 DC vd1_val
Vac d1 d10 AC 1

.DC Vd1 LIN 1 vd1_val vd1_val SWEEP DATA=datanm

.AC LIN 1 10k 10k SWEEP DATA=datanm
.measure ac real_v param = 'VR(d1)' 
.measure ac imag_v param = 'VI(d1)' 
.measure ac real_i param = 'IR(Vac)'
.measure ac imag_i param = 'II(Vac)'
.measure dc Idc1 find i(Vd1) when v(d1)=vd1_val
.measure dc Idc0 find i(Vd0) when v(d1)=vd1_val

.DATA datanm
+ vd0_val vd1_val
+ 0.0 0.0
+ 0.0 0.042105263157894736
+ 0.0 0.08421052631578947
+ 0.0 0.12631578947368421
+ 0.0 0.16842105263157894
+ 0.0 0.21052631578947367
+ 0.0 0.25263157894736843
+ 0.0 0.29473684210526313
+ 0.0 0.3368421052631579
+ 0.0 0.37894736842105264
+ 0.0 0.42105263157894735
+ 0.0 0.4631578947368421
+ 0.0 0.5052631578947369
+ 0.0 0.5473684210526316
+ 0.0 0.5894736842105263
+ 0.0 0.631578947368421
+ 0.0 0.6736842105263158
+ 0.0 0.7157894736842105
+ 0.0 0.7578947368421053
+ 0.0 0.8
+ 0.042105263157894736 0.0
+ 0.042105263157894736 0.042105263157894736
+ 0.042105263157894736 0.08421052631578947
+ 0.042105263157894736 0.12631578947368421
+ 0.042105263157894736 0.16842105263157894
+ 0.042105263157894736 0.21052631578947367
+ 0.042105263157894736 0.25263157894736843
+ 0.042105263157894736 0.29473684210526313
+ 0.042105263157894736 0.3368421052631579
+ 0.042105263157894736 0.37894736842105264
+ 0.042105263157894736 0.42105263157894735
+ 0.042105263157894736 0.4631578947368421
+ 0.042105263157894736 0.5052631578947369
+ 0.042105263157894736 0.5473684210526316
+ 0.042105263157894736 0.5894736842105263
+ 0.042105263157894736 0.631578947368421
+ 0.042105263157894736 0.6736842105263158
+ 0.042105263157894736 0.7157894736842105
+ 0.042105263157894736 0.7578947368421053
+ 0.042105263157894736 0.8
+ 0.08421052631578947 0.0
+ 0.08421052631578947 0.042105263157894736
+ 0.08421052631578947 0.08421052631578947
+ 0.08421052631578947 0.12631578947368421
+ 0.08421052631578947 0.16842105263157894
+ 0.08421052631578947 0.21052631578947367
+ 0.08421052631578947 0.25263157894736843
+ 0.08421052631578947 0.29473684210526313
+ 0.08421052631578947 0.3368421052631579
+ 0.08421052631578947 0.37894736842105264
+ 0.08421052631578947 0.42105263157894735
+ 0.08421052631578947 0.4631578947368421
+ 0.08421052631578947 0.5052631578947369
+ 0.08421052631578947 0.5473684210526316
+ 0.08421052631578947 0.5894736842105263
+ 0.08421052631578947 0.631578947368421
+ 0.08421052631578947 0.6736842105263158
+ 0.08421052631578947 0.7157894736842105
+ 0.08421052631578947 0.7578947368421053
+ 0.08421052631578947 0.8
+ 0.12631578947368421 0.0
+ 0.12631578947368421 0.042105263157894736
+ 0.12631578947368421 0.08421052631578947
+ 0.12631578947368421 0.12631578947368421
+ 0.12631578947368421 0.16842105263157894
+ 0.12631578947368421 0.21052631578947367
+ 0.12631578947368421 0.25263157894736843
+ 0.12631578947368421 0.29473684210526313
+ 0.12631578947368421 0.3368421052631579
+ 0.12631578947368421 0.37894736842105264
+ 0.12631578947368421 0.42105263157894735
+ 0.12631578947368421 0.4631578947368421
+ 0.12631578947368421 0.5052631578947369
+ 0.12631578947368421 0.5473684210526316
+ 0.12631578947368421 0.5894736842105263
+ 0.12631578947368421 0.631578947368421
+ 0.12631578947368421 0.6736842105263158
+ 0.12631578947368421 0.7157894736842105
+ 0.12631578947368421 0.7578947368421053
+ 0.12631578947368421 0.8
+ 0.16842105263157894 0.0
+ 0.16842105263157894 0.042105263157894736
+ 0.16842105263157894 0.08421052631578947
+ 0.16842105263157894 0.12631578947368421
+ 0.16842105263157894 0.16842105263157894
+ 0.16842105263157894 0.21052631578947367
+ 0.16842105263157894 0.25263157894736843
+ 0.16842105263157894 0.29473684210526313
+ 0.16842105263157894 0.3368421052631579
+ 0.16842105263157894 0.37894736842105264
+ 0.16842105263157894 0.42105263157894735
+ 0.16842105263157894 0.4631578947368421
+ 0.16842105263157894 0.5052631578947369
+ 0.16842105263157894 0.5473684210526316
+ 0.16842105263157894 0.5894736842105263
+ 0.16842105263157894 0.631578947368421
+ 0.16842105263157894 0.6736842105263158
+ 0.16842105263157894 0.7157894736842105
+ 0.16842105263157894 0.7578947368421053
+ 0.16842105263157894 0.8
+ 0.21052631578947367 0.0
+ 0.21052631578947367 0.042105263157894736
+ 0.21052631578947367 0.08421052631578947
+ 0.21052631578947367 0.12631578947368421
+ 0.21052631578947367 0.16842105263157894
+ 0.21052631578947367 0.21052631578947367
+ 0.21052631578947367 0.25263157894736843
+ 0.21052631578947367 0.29473684210526313
+ 0.21052631578947367 0.3368421052631579
+ 0.21052631578947367 0.37894736842105264
+ 0.21052631578947367 0.42105263157894735
+ 0.21052631578947367 0.4631578947368421
+ 0.21052631578947367 0.5052631578947369
+ 0.21052631578947367 0.5473684210526316
+ 0.21052631578947367 0.5894736842105263
+ 0.21052631578947367 0.631578947368421
+ 0.21052631578947367 0.6736842105263158
+ 0.21052631578947367 0.7157894736842105
+ 0.21052631578947367 0.7578947368421053
+ 0.21052631578947367 0.8
+ 0.25263157894736843 0.0
+ 0.25263157894736843 0.042105263157894736
+ 0.25263157894736843 0.08421052631578947
+ 0.25263157894736843 0.12631578947368421
+ 0.25263157894736843 0.16842105263157894
+ 0.25263157894736843 0.21052631578947367
+ 0.25263157894736843 0.25263157894736843
+ 0.25263157894736843 0.29473684210526313
+ 0.25263157894736843 0.3368421052631579
+ 0.25263157894736843 0.37894736842105264
+ 0.25263157894736843 0.42105263157894735
+ 0.25263157894736843 0.4631578947368421
+ 0.25263157894736843 0.5052631578947369
+ 0.25263157894736843 0.5473684210526316
+ 0.25263157894736843 0.5894736842105263
+ 0.25263157894736843 0.631578947368421
+ 0.25263157894736843 0.6736842105263158
+ 0.25263157894736843 0.7157894736842105
+ 0.25263157894736843 0.7578947368421053
+ 0.25263157894736843 0.8
+ 0.29473684210526313 0.0
+ 0.29473684210526313 0.042105263157894736
+ 0.29473684210526313 0.08421052631578947
+ 0.29473684210526313 0.12631578947368421
+ 0.29473684210526313 0.16842105263157894
+ 0.29473684210526313 0.21052631578947367
+ 0.29473684210526313 0.25263157894736843
+ 0.29473684210526313 0.29473684210526313
+ 0.29473684210526313 0.3368421052631579
+ 0.29473684210526313 0.37894736842105264
+ 0.29473684210526313 0.42105263157894735
+ 0.29473684210526313 0.4631578947368421
+ 0.29473684210526313 0.5052631578947369
+ 0.29473684210526313 0.5473684210526316
+ 0.29473684210526313 0.5894736842105263
+ 0.29473684210526313 0.631578947368421
+ 0.29473684210526313 0.6736842105263158
+ 0.29473684210526313 0.7157894736842105
+ 0.29473684210526313 0.7578947368421053
+ 0.29473684210526313 0.8
+ 0.3368421052631579 0.0
+ 0.3368421052631579 0.042105263157894736
+ 0.3368421052631579 0.08421052631578947
+ 0.3368421052631579 0.12631578947368421
+ 0.3368421052631579 0.16842105263157894
+ 0.3368421052631579 0.21052631578947367
+ 0.3368421052631579 0.25263157894736843
+ 0.3368421052631579 0.29473684210526313
+ 0.3368421052631579 0.3368421052631579
+ 0.3368421052631579 0.37894736842105264
+ 0.3368421052631579 0.42105263157894735
+ 0.3368421052631579 0.4631578947368421
+ 0.3368421052631579 0.5052631578947369
+ 0.3368421052631579 0.5473684210526316
+ 0.3368421052631579 0.5894736842105263
+ 0.3368421052631579 0.631578947368421
+ 0.3368421052631579 0.6736842105263158
+ 0.3368421052631579 0.7157894736842105
+ 0.3368421052631579 0.7578947368421053
+ 0.3368421052631579 0.8
+ 0.37894736842105264 0.0
+ 0.37894736842105264 0.042105263157894736
+ 0.37894736842105264 0.08421052631578947
+ 0.37894736842105264 0.12631578947368421
+ 0.37894736842105264 0.16842105263157894
+ 0.37894736842105264 0.21052631578947367
+ 0.37894736842105264 0.25263157894736843
+ 0.37894736842105264 0.29473684210526313
+ 0.37894736842105264 0.3368421052631579
+ 0.37894736842105264 0.37894736842105264
+ 0.37894736842105264 0.42105263157894735
+ 0.37894736842105264 0.4631578947368421
+ 0.37894736842105264 0.5052631578947369
+ 0.37894736842105264 0.5473684210526316
+ 0.37894736842105264 0.5894736842105263
+ 0.37894736842105264 0.631578947368421
+ 0.37894736842105264 0.6736842105263158
+ 0.37894736842105264 0.7157894736842105
+ 0.37894736842105264 0.7578947368421053
+ 0.37894736842105264 0.8
+ 0.42105263157894735 0.0
+ 0.42105263157894735 0.042105263157894736
+ 0.42105263157894735 0.08421052631578947
+ 0.42105263157894735 0.12631578947368421
+ 0.42105263157894735 0.16842105263157894
+ 0.42105263157894735 0.21052631578947367
+ 0.42105263157894735 0.25263157894736843
+ 0.42105263157894735 0.29473684210526313
+ 0.42105263157894735 0.3368421052631579
+ 0.42105263157894735 0.37894736842105264
+ 0.42105263157894735 0.42105263157894735
+ 0.42105263157894735 0.4631578947368421
+ 0.42105263157894735 0.5052631578947369
+ 0.42105263157894735 0.5473684210526316
+ 0.42105263157894735 0.5894736842105263
+ 0.42105263157894735 0.631578947368421
+ 0.42105263157894735 0.6736842105263158
+ 0.42105263157894735 0.7157894736842105
+ 0.42105263157894735 0.7578947368421053
+ 0.42105263157894735 0.8
+ 0.4631578947368421 0.0
+ 0.4631578947368421 0.042105263157894736
+ 0.4631578947368421 0.08421052631578947
+ 0.4631578947368421 0.12631578947368421
+ 0.4631578947368421 0.16842105263157894
+ 0.4631578947368421 0.21052631578947367
+ 0.4631578947368421 0.25263157894736843
+ 0.4631578947368421 0.29473684210526313
+ 0.4631578947368421 0.3368421052631579
+ 0.4631578947368421 0.37894736842105264
+ 0.4631578947368421 0.42105263157894735
+ 0.4631578947368421 0.4631578947368421
+ 0.4631578947368421 0.5052631578947369
+ 0.4631578947368421 0.5473684210526316
+ 0.4631578947368421 0.5894736842105263
+ 0.4631578947368421 0.631578947368421
+ 0.4631578947368421 0.6736842105263158
+ 0.4631578947368421 0.7157894736842105
+ 0.4631578947368421 0.7578947368421053
+ 0.4631578947368421 0.8
+ 0.5052631578947369 0.0
+ 0.5052631578947369 0.042105263157894736
+ 0.5052631578947369 0.08421052631578947
+ 0.5052631578947369 0.12631578947368421
+ 0.5052631578947369 0.16842105263157894
+ 0.5052631578947369 0.21052631578947367
+ 0.5052631578947369 0.25263157894736843
+ 0.5052631578947369 0.29473684210526313
+ 0.5052631578947369 0.3368421052631579
+ 0.5052631578947369 0.37894736842105264
+ 0.5052631578947369 0.42105263157894735
+ 0.5052631578947369 0.4631578947368421
+ 0.5052631578947369 0.5052631578947369
+ 0.5052631578947369 0.5473684210526316
+ 0.5052631578947369 0.5894736842105263
+ 0.5052631578947369 0.631578947368421
+ 0.5052631578947369 0.6736842105263158
+ 0.5052631578947369 0.7157894736842105
+ 0.5052631578947369 0.7578947368421053
+ 0.5052631578947369 0.8
+ 0.5473684210526316 0.0
+ 0.5473684210526316 0.042105263157894736
+ 0.5473684210526316 0.08421052631578947
+ 0.5473684210526316 0.12631578947368421
+ 0.5473684210526316 0.16842105263157894
+ 0.5473684210526316 0.21052631578947367
+ 0.5473684210526316 0.25263157894736843
+ 0.5473684210526316 0.29473684210526313
+ 0.5473684210526316 0.3368421052631579
+ 0.5473684210526316 0.37894736842105264
+ 0.5473684210526316 0.42105263157894735
+ 0.5473684210526316 0.4631578947368421
+ 0.5473684210526316 0.5052631578947369
+ 0.5473684210526316 0.5473684210526316
+ 0.5473684210526316 0.5894736842105263
+ 0.5473684210526316 0.631578947368421
+ 0.5473684210526316 0.6736842105263158
+ 0.5473684210526316 0.7157894736842105
+ 0.5473684210526316 0.7578947368421053
+ 0.5473684210526316 0.8
+ 0.5894736842105263 0.0
+ 0.5894736842105263 0.042105263157894736
+ 0.5894736842105263 0.08421052631578947
+ 0.5894736842105263 0.12631578947368421
+ 0.5894736842105263 0.16842105263157894
+ 0.5894736842105263 0.21052631578947367
+ 0.5894736842105263 0.25263157894736843
+ 0.5894736842105263 0.29473684210526313
+ 0.5894736842105263 0.3368421052631579
+ 0.5894736842105263 0.37894736842105264
+ 0.5894736842105263 0.42105263157894735
+ 0.5894736842105263 0.4631578947368421
+ 0.5894736842105263 0.5052631578947369
+ 0.5894736842105263 0.5473684210526316
+ 0.5894736842105263 0.5894736842105263
+ 0.5894736842105263 0.631578947368421
+ 0.5894736842105263 0.6736842105263158
+ 0.5894736842105263 0.7157894736842105
+ 0.5894736842105263 0.7578947368421053
+ 0.5894736842105263 0.8
+ 0.631578947368421 0.0
+ 0.631578947368421 0.042105263157894736
+ 0.631578947368421 0.08421052631578947
+ 0.631578947368421 0.12631578947368421
+ 0.631578947368421 0.16842105263157894
+ 0.631578947368421 0.21052631578947367
+ 0.631578947368421 0.25263157894736843
+ 0.631578947368421 0.29473684210526313
+ 0.631578947368421 0.3368421052631579
+ 0.631578947368421 0.37894736842105264
+ 0.631578947368421 0.42105263157894735
+ 0.631578947368421 0.4631578947368421
+ 0.631578947368421 0.5052631578947369
+ 0.631578947368421 0.5473684210526316
+ 0.631578947368421 0.5894736842105263
+ 0.631578947368421 0.631578947368421
+ 0.631578947368421 0.6736842105263158
+ 0.631578947368421 0.7157894736842105
+ 0.631578947368421 0.7578947368421053
+ 0.631578947368421 0.8
+ 0.6736842105263158 0.0
+ 0.6736842105263158 0.042105263157894736
+ 0.6736842105263158 0.08421052631578947
+ 0.6736842105263158 0.12631578947368421
+ 0.6736842105263158 0.16842105263157894
+ 0.6736842105263158 0.21052631578947367
+ 0.6736842105263158 0.25263157894736843
+ 0.6736842105263158 0.29473684210526313
+ 0.6736842105263158 0.3368421052631579
+ 0.6736842105263158 0.37894736842105264
+ 0.6736842105263158 0.42105263157894735
+ 0.6736842105263158 0.4631578947368421
+ 0.6736842105263158 0.5052631578947369
+ 0.6736842105263158 0.5473684210526316
+ 0.6736842105263158 0.5894736842105263
+ 0.6736842105263158 0.631578947368421
+ 0.6736842105263158 0.6736842105263158
+ 0.6736842105263158 0.7157894736842105
+ 0.6736842105263158 0.7578947368421053
+ 0.6736842105263158 0.8
+ 0.7157894736842105 0.0
+ 0.7157894736842105 0.042105263157894736
+ 0.7157894736842105 0.08421052631578947
+ 0.7157894736842105 0.12631578947368421
+ 0.7157894736842105 0.16842105263157894
+ 0.7157894736842105 0.21052631578947367
+ 0.7157894736842105 0.25263157894736843
+ 0.7157894736842105 0.29473684210526313
+ 0.7157894736842105 0.3368421052631579
+ 0.7157894736842105 0.37894736842105264
+ 0.7157894736842105 0.42105263157894735
+ 0.7157894736842105 0.4631578947368421
+ 0.7157894736842105 0.5052631578947369
+ 0.7157894736842105 0.5473684210526316
+ 0.7157894736842105 0.5894736842105263
+ 0.7157894736842105 0.631578947368421
+ 0.7157894736842105 0.6736842105263158
+ 0.7157894736842105 0.7157894736842105
+ 0.7157894736842105 0.7578947368421053
+ 0.7157894736842105 0.8
+ 0.7578947368421053 0.0
+ 0.7578947368421053 0.042105263157894736
+ 0.7578947368421053 0.08421052631578947
+ 0.7578947368421053 0.12631578947368421
+ 0.7578947368421053 0.16842105263157894
+ 0.7578947368421053 0.21052631578947367
+ 0.7578947368421053 0.25263157894736843
+ 0.7578947368421053 0.29473684210526313
+ 0.7578947368421053 0.3368421052631579
+ 0.7578947368421053 0.37894736842105264
+ 0.7578947368421053 0.42105263157894735
+ 0.7578947368421053 0.4631578947368421
+ 0.7578947368421053 0.5052631578947369
+ 0.7578947368421053 0.5473684210526316
+ 0.7578947368421053 0.5894736842105263
+ 0.7578947368421053 0.631578947368421
+ 0.7578947368421053 0.6736842105263158
+ 0.7578947368421053 0.7157894736842105
+ 0.7578947368421053 0.7578947368421053
+ 0.7578947368421053 0.8
+ 0.8 0.0
+ 0.8 0.042105263157894736
+ 0.8 0.08421052631578947
+ 0.8 0.12631578947368421
+ 0.8 0.16842105263157894
+ 0.8 0.21052631578947367
+ 0.8 0.25263157894736843
+ 0.8 0.29473684210526313
+ 0.8 0.3368421052631579
+ 0.8 0.37894736842105264
+ 0.8 0.42105263157894735
+ 0.8 0.4631578947368421
+ 0.8 0.5052631578947369
+ 0.8 0.5473684210526316
+ 0.8 0.5894736842105263
+ 0.8 0.631578947368421
+ 0.8 0.6736842105263158
+ 0.8 0.7157894736842105
+ 0.8 0.7578947368421053
+ 0.8 0.8
.ENDDATA

.end
