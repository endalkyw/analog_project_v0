.subckt nmos_cm_1 d0 d1 s 
* Net:s ----------------
R1 s s:27 3.108
R2 s s:26 0.42
R3 s s:19 1.092
R4 s s:2 4.368
R5 s:2 s:31 3.108
R6 s:2 MN0@2:s 14
R7 s:2 s:30 0.42
R8 s:2 MN0@2:s 14
R9 s:2 s:1 4.368
R10 s:2 MN0@2:s 14
R11 s:2 s:6 3.724
R12 s:2 MN0@2:s 14
R13 s:6 s:0 18.984
R14 s:6 s:3 0.644
R15 s:3 s:35 3.108
R16 s:3 MN1@2:s 14
R17 s:3 s:34 0.42
R18 s:3 MN1@2:s 14
R19 s:3 s:4 4.368
R20 s:3 MN1@2:s 14
R21 s:4 s:39 3.108
R22 s:4 MN0@4:s 14
R23 s:4 s:38 0.42
R24 s:4 MN0@4:s 14
R25 s:4 s:5 4.368
R26 s:4 MN0@4:s 14
R27 s:5 s:43 3.108
R28 s:5 MN1@4:s 14
R29 s:5 s:42 0.42
R30 s:5 MN1@4:s 14
R31 s:5 s:20 1.092
R32 s:5 MN1@4:s 14
R33 s:42 s:17 1.708
R34 s:42 MN1@4:s 14
R35 s:43 s:44 3.528
R36 s:43 MN1@4:s 14
R37 s:44 s:45 3.528
R38 s:44 MN1@4:s 14
R39 s:45 s:18 1.428
R40 s:45 MN1@4:s 14
R41 s:38 s:15 1.708
R42 s:38 MN0@4:s 14
R43 s:39 s:40 3.528
R44 s:39 MN0@4:s 14
R45 s:40 s:41 3.528
R46 s:40 MN0@4:s 14
R47 s:41 s:16 1.428
R48 s:41 MN0@4:s 14
R49 s:34 s:13 1.708
R50 s:34 MN1@2:s 14
R51 s:35 s:36 3.528
R52 s:35 MN1@2:s 14
R53 s:36 s:37 3.528
R54 s:36 MN1@2:s 14
R55 s:37 s:14 1.428
R56 s:37 MN1@2:s 14
R57 s:0 s:21 1.176
R58 s:0 MN0:b 14
R59 s:0 s:23 1.12
R60 s:0 MN0:b 14
R61 s:0 s:24 2.408
R62 s:0 MN0:b 14
R63 s:24 s:25 3.528
R64 s:24 MN0:b 14
R65 s:25 s:8 1.59
R66 s:25 MN0:b 14
R67 s:23 s:22 3.528
R68 s:23 MN0:b 14
R69 s:22 s:7 1.59
R70 s:22 MN0:b 14
R71 s:1 s:27 3.108
R72 s:1 MN0:s 14
R73 s:1 s:26 0.42
R74 s:1 MN0:s 14
R75 s:1 s:19 1.092
R76 s:1 MN0:s 14
R77 s:26 s:9 1.708
R78 s:26 MN0:s 14
R79 s:27 s:28 3.528
R80 s:27 MN0:s 14
R81 s:28 s:29 3.528
R82 s:28 MN0:s 14
R83 s:29 s:10 1.428
R84 s:29 MN0:s 14
R85 s:30 s:11 1.708
R86 s:30 MN0@2:s 14
R87 s:31 s:32 3.528
R88 s:31 MN0@2:s 14
R89 s:32 s:33 3.528
R90 s:32 MN0@2:s 14
R91 s:33 s:12 1.428
R92 s:33 MN0@2:s 14
R93 MN0:b MN0@2:b 0.01
R94 MN0@2:b MN1:b 0.01
R95 MN1:b MN1@2:b 0.01
R96 MN1@2:b MN0@3:b 0.01
R97 MN0@3:b MN0@4:b 0.01
R98 MN0@4:b MN1@3:b 0.01
R99 MN1@3:b MN1@4:b 0.01
R100 MN0@2:s MN1:s 0.01
R101 MN1@2:s MN0@3:s 0.01
R102 MN0@4:s MN1@3:s 0.01
C1 s:2 0 2.331e-14
C2 s:2 0 3.1500000000000003e-15
C3 s:2 0 3.2760000000000004e-14
C4 s:2 0 2.793e-14
C5 s:6 0 1.4238e-13
C6 s:6 0 4.83e-15
C7 s:3 0 2.331e-14
C8 s:3 0 3.1500000000000003e-15
C9 s:3 0 3.2760000000000004e-14
C10 s:4 0 2.331e-14
C11 s:4 0 3.1500000000000003e-15
C12 s:4 0 3.2760000000000004e-14
C13 s:5 0 2.331e-14
C14 s:5 0 3.1500000000000003e-15
C15 s:5 0 8.190000000000001e-15
C16 s:42 0 1.2810000000000001e-14
C17 s:43 0 2.6460000000000002e-14
C18 s:44 0 2.6460000000000002e-14
C19 s:45 0 1.0710000000000001e-14
C20 s:38 0 1.2810000000000001e-14
C21 s:39 0 2.6460000000000002e-14
C22 s:40 0 2.6460000000000002e-14
C23 s:41 0 1.0710000000000001e-14
C24 s:34 0 1.2810000000000001e-14
C25 s:35 0 2.6460000000000002e-14
C26 s:36 0 2.6460000000000002e-14
C27 s:37 0 1.0710000000000001e-14
C28 s:0 0 8.82e-15
C29 s:0 0 8.400000000000001e-15
C30 s:0 0 1.806e-14
C31 s:24 0 2.6460000000000002e-14
C32 s:25 0 1.1928000000000016e-14
C33 s:23 0 2.6460000000000002e-14
C34 s:22 0 1.1928000000000003e-14
C35 s:1 0 2.331e-14
C36 s:1 0 3.1500000000000003e-15
C37 s:1 0 8.190000000000001e-15
C38 s:26 0 1.2810000000000001e-14
C39 s:27 0 2.6460000000000002e-14
C40 s:28 0 2.6460000000000002e-14
C41 s:29 0 1.0710000000000001e-14
C42 s:30 0 1.2810000000000001e-14
C43 s:31 0 2.6460000000000002e-14
C44 s:32 0 2.6460000000000002e-14
C45 s:33 0 1.0710000000000001e-14

* Net:d0 ----------------
R103 d0 d0:6 0.98
R104 d0 d0:2 0.728
R105 d0:6 d0:7 3.528
R106 d0:6 MN0:d 14
R107 d0:7 d0:8 3.528
R108 d0:7 MN0:d 14
R109 d0:8 d0:9 3.528
R110 d0:8 MN0:d 14
R111 d0:9 d0:0 3.696
R112 d0:9 MN0:d 14
R113 d0:0 d0:14 0.294
R114 d0:0 MN0:g 342
R115 d0:0 MN0@2:g 342
R116 d0:0 MN1:g 342
R117 d0:0 MN1@2:g 342
R118 d0:0 MN0@3:g 342
R119 d0:0 MN0@4:g 342
R120 d0:0 MN1@3:g 342
R121 d0:0 MN1@4:g 342
R122 d0:0 d0:15 3.234
R123 d0:0 MN0:g 342
R124 d0:0 MN0@2:g 342
R125 d0:0 MN1:g 342
R126 d0:0 MN1@2:g 342
R127 d0:0 MN0@3:g 342
R128 d0:0 MN0@4:g 342
R129 d0:0 MN1@3:g 342
R130 d0:0 MN1@4:g 342
R131 d0:15 d0:16 3.528
R132 d0:15 MN0:g 342
R133 d0:15 MN0@2:g 342
R134 d0:15 MN1:g 342
R135 d0:15 MN1@2:g 342
R136 d0:15 MN0@3:g 342
R137 d0:15 MN0@4:g 342
R138 d0:15 MN1@3:g 342
R139 d0:15 MN1@4:g 342
R140 d0:16 d0:1 1.974
R141 d0:16 MN0:g 342
R142 d0:16 MN0@2:g 342
R143 d0:16 MN1:g 342
R144 d0:16 MN1@2:g 342
R145 d0:16 MN0@3:g 342
R146 d0:16 MN0@4:g 342
R147 d0:16 MN1@3:g 342
R148 d0:16 MN1@4:g 342
R149 d0:1 d0:13 3.696
R150 d0:1 MN0:g 342
R151 d0:1 MN0@2:g 342
R152 d0:1 MN1:g 342
R153 d0:1 MN1@2:g 342
R154 d0:1 MN0@3:g 342
R155 d0:1 MN0@4:g 342
R156 d0:1 MN1@3:g 342
R157 d0:1 MN1@4:g 342
R158 d0:1 d0:17 1.554
R159 d0:1 MN0:g 342
R160 d0:1 MN0@2:g 342
R161 d0:1 MN1:g 342
R162 d0:1 MN1@2:g 342
R163 d0:1 MN0@3:g 342
R164 d0:1 MN0@4:g 342
R165 d0:1 MN1@3:g 342
R166 d0:1 MN1@4:g 342
R167 d0:17 d0:18 3.528
R168 d0:17 MN0:g 342
R169 d0:17 MN0@2:g 342
R170 d0:17 MN1:g 342
R171 d0:17 MN1@2:g 342
R172 d0:17 MN0@3:g 342
R173 d0:17 MN0@4:g 342
R174 d0:17 MN1@3:g 342
R175 d0:17 MN1@4:g 342
R176 d0:18 d0:5 2.562
R177 d0:18 MN0:g 342
R178 d0:18 MN0@2:g 342
R179 d0:18 MN1:g 342
R180 d0:18 MN1@2:g 342
R181 d0:18 MN0@3:g 342
R182 d0:18 MN0@4:g 342
R183 d0:18 MN1@3:g 342
R184 d0:18 MN1@4:g 342
R185 d0:13 d0:12 3.528
R186 d0:13 MN0@3:d 14
R187 d0:12 d0:11 3.528
R188 d0:12 MN0@3:d 14
R189 d0:11 d0:10 3.528
R190 d0:11 MN0@3:d 14
R191 d0:10 d0:3 1.708
R192 d0:10 MN0@3:d 14
R193 d0:14 d0:4 2.982
R194 d0:14 MN0:g 342
R195 d0:14 MN0@2:g 342
R196 d0:14 MN1:g 342
R197 d0:14 MN1@2:g 342
R198 d0:14 MN0@3:g 342
R199 d0:14 MN0@4:g 342
R200 d0:14 MN1@3:g 342
R201 d0:14 MN1@4:g 342
R202 MN0:d MN0@2:d 0.01
R203 MN0@3:d MN0@4:d 0.01
C46 d0:6 0 2.6460000000000002e-14
C47 d0:7 0 2.6460000000000002e-14
C48 d0:8 0 2.6460000000000002e-14
C49 d0:9 0 2.772e-14
C50 d0:0 0 2.205e-15
C51 d0:0 0 2.4255e-14
C52 d0:15 0 2.6460000000000002e-14
C53 d0:16 0 1.4805e-14
C54 d0:1 0 2.772e-14
C55 d0:1 0 1.1655e-14
C56 d0:17 0 2.6460000000000002e-14
C57 d0:18 0 1.9215e-14
C58 d0:13 0 2.6460000000000002e-14
C59 d0:12 0 2.6460000000000002e-14
C60 d0:11 0 2.6460000000000002e-14
C61 d0:10 0 1.2810000000000001e-14
C62 d0:14 0 2.2365e-14


* Net:d1 ----------------
R204 d1 d1:8 2.66
R205 d1 d1:2 0.588
R206 d1 d1:6 0.728
R207 d1 d1:1 8.736
R208 d1:1 d1:12 2.66
R209 d1:1 d1:4 0.588
R210 d1:1 d1:0 8.736
R211 d1:1 d1:7 0.728
R212 d1:0 d1:8 2.66
R213 d1:0 d1:2 0.588
R214 d1:0 d1:6 0.728
R215 d1:8 d1:9 3.528
R216 d1:8 MN1:d 14
R217 d1:9 d1:10 3.528
R218 d1:9 MN1:d 14
R219 d1:10 d1:11 3.528
R220 d1:10 MN1:d 14
R221 d1:11 d1:3 1.428
R222 d1:11 MN1:d 14
R223 d1:12 d1:13 3.528
R224 d1:12 MN1@3:d 14
R225 d1:13 d1:14 3.528
R226 d1:13 MN1@3:d 14
R227 d1:14 d1:15 3.528
R228 d1:14 MN1@3:d 14
R229 d1:15 d1:5 1.428
R230 d1:15 MN1@3:d 14
R231 MN1:d MN1@2:d 0.01
R232 MN1@3:d MN1@4:d 0.01
C63 d1:1 0 1.995e-14
C64 d1:1 0 4.41e-15
C65 d1:1 0 6.552000000000001e-14
C66 d1:1 0 5.46e-15
C67 d1:0 0 1.995e-14
C68 d1:0 0 4.41e-15
C69 d1:0 0 5.46e-15
C70 d1:8 0 2.6460000000000002e-14
C71 d1:9 0 2.6460000000000002e-14
C72 d1:10 0 2.6460000000000002e-14
C73 d1:11 0 1.0710000000000001e-14
C74 d1:12 0 2.6460000000000002e-14
C75 d1:13 0 2.6460000000000002e-14
C76 d1:14 0 2.6460000000000002e-14
C77 d1:15 0 1.0710000000000001e-14

XXMN0 MN0:d MN0:g MN0:s MN0:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10 nf=1
+ plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1 par=1
+ dtemp=0 l_shape=0 l_shape_s=0 asej=5.94e-15 adej=2.97e-15 psej=1.19e-06
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=6.17e-07
+ lle_sb=7.1e-08 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.383e-06 lle_rxrxb=1.929e-06 lle_rxrxs=1e-06 lle_rxrxn=6.42197e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=8.19e-07 lle_ctse=8.19e-07
+ lle_ctnw=2.73e-07 lle_ctsw=2.73e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.252 $Y=0.127
XXMN0@2 MN0@4:d MN0@4:g MN0@4:s MN0@4:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=2.97e-15 psej=5.4e-07
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=5.39e-07
+ lle_sb=1.49e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.461e-06 lle_rxrxb=1.851e-06 lle_rxrxs=1e-06 lle_rxrxn=3.19671e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=7.41e-07 lle_ctse=7.41e-07
+ lle_ctnw=3.51e-07 lle_ctsw=3.51e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.33 $Y=0.127
XXMN1 MN1:d MN1:g MN1:s MN1:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10 nf=1
+ plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1 par=1
+ dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=2.97e-15 psej=5.4e-07
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=4.61e-07
+ lle_sb=2.27e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.539e-06 lle_rxrxb=1.773e-06 lle_rxrxs=1e-06 lle_rxrxn=2.34e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=6.63e-07 lle_ctse=6.63e-07
+ lle_ctnw=4.29e-07 lle_ctsw=4.29e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.408 $Y=0.127
XXMN1@2 MN1@4:d MN1@4:g MN1@4:s MN1@4:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=2.97e-15 psej=5.4e-07
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=3.83e-07
+ lle_sb=3.05e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.617e-06 lle_rxrxb=1.695e-06 lle_rxrxs=1e-06 lle_rxrxn=2.34e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=5.85e-07 lle_ctse=5.85e-07
+ lle_ctnw=5.07e-07 lle_ctsw=5.07e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.486 $Y=0.127
XXMN0@3 MN0@3:d MN0@3:g MN0@3:s MN0@3:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=2.97e-15 psej=5.4e-07
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=3.05e-07
+ lle_sb=3.83e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.695e-06 lle_rxrxb=1.617e-06 lle_rxrxs=1e-06 lle_rxrxn=2.34e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=5.07e-07 lle_ctse=5.07e-07
+ lle_ctnw=5.85e-07 lle_ctsw=5.85e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.564 $Y=0.127
XXMN0@4 MN0@2:d MN0@2:g MN0@2:s MN0@2:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=2.97e-15 psej=5.4e-07
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=2.27e-07
+ lle_sb=4.61e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.773e-06 lle_rxrxb=1.539e-06 lle_rxrxs=1e-06 lle_rxrxn=2.34e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=4.29e-07 lle_ctse=4.29e-07
+ lle_ctnw=6.63e-07 lle_ctsw=6.63e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.642 $Y=0.127
XXMN1@3 MN1@3:d MN1@3:g MN1@3:s MN1@3:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=2.97e-15 psej=5.4e-07
+ pdej=5.4e-07 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=1.49e-07
+ lle_sb=5.39e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.851e-06 lle_rxrxb=1.461e-06 lle_rxrxs=1e-06 lle_rxrxn=3.19671e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=3.51e-07 lle_ctse=3.51e-07
+ lle_ctnw=7.41e-07 lle_ctsw=7.41e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.72 $Y=0.127
XXMN1@4 MN1@2:d MN1@2:g MN1@2:s MN1@2:b nfet l=1.4e-08 fpitch=4.8e-08 nfin=10
+ nf=1 plorient=0 p_la=0 ngcon=1 cpp=7.8e-08 analog=-1 nf_pex=4 par_nf=4 m=1
+ par=1 dtemp=0 l_shape=0 l_shape_s=0 asej=2.97e-15 adej=5.94e-15 psej=5.4e-07
+ pdej=1.19e-06 sca=3.65883 scb=0.00013005 scc=4.86669e-09 lle_sa=7.1e-08
+ lle_sb=6.17e-07 lle_nwa=2e-06 lle_nwb=2e-06 lle_nws=2e-06 lle_nwn=2e-06
+ lle_rxrxa=1.929e-06 lle_rxrxb=1.383e-06 lle_rxrxs=1e-06 lle_rxrxn=6.42197e-07
+ lle_pcrxs=5.5e-08 lle_pcrxn=1.07e-07 lle_ctne=2.73e-07 lle_ctse=2.73e-07
+ lle_ctnw=8.19e-07 lle_ctsw=8.19e-07 lle_sctne=0 lle_sctnw=0 lle_sctse=0
+ lle_sctsw=0 ptwell=0 pre_layout_local=0 pre_layout_local_rd=0
+ pre_layout_local_rs=0 pre_layout_local_rg=0 $X=0.798 $Y=0.127


.ends nmos_cm_1
